LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE work.kasumi_pack.ALL;

ENTITY kasumi_tb IS END kasumi_tb;

ARCHITECTURE test OF kasumi_tb IS
	SIGNAL pt:    u64;
	SIGNAL kt:    u128;
	SIGNAL clk:   std_logic;
	SIGNAL nrst:  std_logic;
	SIGNAL ct:    u64;
BEGIN
	dut: ENTITY work.kasumi PORT MAP(
		pt, kt, clk, nrst, ct
	);
	
	PROCESS
	BEGIN
		pt   <= "0000000000000000000000000000000000000000000000000000000000000000";
		kt   <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
		clk  <= '0';
		nrst <= '0';
		wait for 10 ns;
		
		pt   <= "0000000000000000000000000000000000000000000000000001000000100110";
		kt   <= "00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000100";
		clk  <= '1';
		nrst <= '1';
		wait for 10 ns;
	END PROCESS;
	
END test;